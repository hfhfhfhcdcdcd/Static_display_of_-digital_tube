module rw_74HC595 (
    input                       DS          ,
    output      reg[13:0]       Q 
);

endmodule